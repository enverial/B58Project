module CleanupDrawings(Clock, Reset, XIn, XOut, YIn, YOut);