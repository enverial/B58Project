module CleanupDrawings(Clock, Reset, State, XOut, YOut);
  // Used to draw black where the character used to be so it doesn't leave an image
